* ======================================================
* Template TB (uses your NETLIST1.cir subckts)
* Works with server.render_tb() placeholders
* ======================================================

.title Uploaded-subckt waveform demo

* --------- Your global models ----------
.MODEL NMOS_GLOBEL NMOS LEVEL=6
.MODEL PMOS_GLOBEL PMOS LEVEL=6

* --------- Your subckts (converted to PARAMS: for clean instantiation) ----------
* NOT gate
.SUBCKT NOT1 OUTPUT INPUT VDD VSS  PARAMS: WP=2u WN=1u L=0.1u M=1
MP0 OUTPUT INPUT VDD VDD PMOS_GLOBEL W={WP} L={L} M={M}
MN0 OUTPUT INPUT VSS VSS NMOS_GLOBEL W={WN} L={L} M={M}
.ENDS NOT1

* 2-input NAND
.SUBCKT NAND2 OUTPUT INPUT1 INPUT2 VDD VSS  PARAMS: WP=2u WN=1u L=0.1u M=1
MP0 OUTPUT INPUT1 VDD VDD PMOS_GLOBEL W={WP} L={L} M={M}
MP1 OUTPUT INPUT2 VDD VDD PMOS_GLOBEL W={WP} L={L} M={M}
MN0 OUTPUT INPUT1 NET1 VSS NMOS_GLOBEL W={WN} L={L} M={M}
MN1 NET1   INPUT2 VSS VSS NMOS_GLOBEL W={WN} L={L} M={M}
.ENDS NAND2

* (Optional) Your higher-level subckt from NETLIST1.cir, kept here if needed
* .SUBCKT NETLIST1 INPUT1 INPUT2 OUTPUT
* XNAND1 NET3 INPUT1 NET2 VDD VSS NAND2 WP=2u WN=1u L=0.1u M=1
* XNAND2 NET3 INPUT2 NET5 VDD VSS NAND2 WP=2u WN=1u L=0.1u M=1
* XNOT1  OUTPUT NET3 VDD VSS NOT1  WP=2u WN=1u L=0.1u M=1
* .ENDS NETLIST1

* --------- Params filled by backend ---------
.param VDD={VDD}
.param TR={TR}
.param TF={TF}
.param PW={PW}
.param PER={PER}
.param CLOAD={CLOAD}
.temp {TEMP}

* --------- Sources ---------
VDD  VDD  0  {VDD}
* /simulate expects ONE driven input → map {A_NODE} to input
VIN  {A_NODE}  0  PULSE(0 {VDD} 0 {TR} {TF} {PW} {PER})

* --------- DUT selection (default: NOT1) ---------
* Single-input flow → NOT1 fits perfectly
XU1  {Y_NODE} {A_NODE} VDD 0  NOT1

* (If you later want NAND2 here, add a second input node and source in code)
* Example (commented):
* VINB  B 0 0
* XU1   {Y_NODE} {A_NODE} B VDD 0 NAND2

* --------- Load & analysis ---------
Cout {Y_NODE}  0  {CLOAD}

.options method=trap reltol=1e-3 abstol=1e-12 vabstol=1e-6 iabstol=1e-12
.options maxord=2

.tran {TSTEP} {TSTOP}
.save time {SAVE_VECTORS}

.control
  set wr_singlescale
  set filetype=ascii
  run
  wrdata {OUT_CSV} time {SAVE_VECTORS}
  * plot v({A_NODE}) v({Y_NODE})
.endc

.end
