* === Uploaded Netlist ===
* Netlist Data

.MODEL NMOS_GLOBEL NMOS LEVEL=6
.MODEL PMOS_GLOBEL PMOS LEVEL=6


.SUBCKT NOT1 OUTPUT INPUT VDD VSS PARAMS: WP=2e-6 WN=1e-6 L=1e-6 M=1
MP0 OUTPUT INPUT VDD VDD PMOS_GLOBEL W=WP L=L M=M
MN0 OUTPUT INPUT VSS VSS NMOS_GLOBEL W=WN L=L M=M
.ENDS

.SUBCKT NAND2 OUTPUT INPUT1 INPUT2 VDD VSS PARAMS: WP=2e-6 WN=1e-6 L=1e-6 M=1
MP0 OUTPUT INPUT1 VDD VDD PMOS_GLOBEL W=WP L=L M=M
MP1 OUTPUT INPUT2 VDD VDD PMOS_GLOBEL W=WP L=L M=M
MN0 OUTPUT INPUT1 NET1 VSS NMOS_GLOBEL W=WN L=L M=M
MN1 NET1   INPUT2 VSS VSS NMOS_GLOBEL W=WN L=L M=M
.ENDS





.SUBCKT NETLIST3 INPUT1 INPUT2 OUTPUT
XNAND1 NET3 INPUT1 NET2 VDD1 VSS1 NAND2 WP=0.000002 WN=0.000001 L=0.000001 M=1
XNAND2 NET3 INPUT2 NET5 VDD2 VSS2 NAND2 WP=0.000002 WN=0.000001 L=0.000001 M=1
XNOT1 OUTPUT NET3 VDD VSS NOT1 WP=0.000002 WN=0.000001 L=0.000001 M=1
XDESIGN1 OUTPUT INPUT1 INPUT2 VDD1 VDD2 VDD VSS1 VSS2 VSS DESIGN1
.ENDS


* === Auto-generated Testbench ===
.options method=trap reltol=1e-3 maxord=2
.temp 25.0

* Sources
VDD VDD 0 1.2
VIN_INPUT2 INPUT2 0 PULSE(0 1.2 0 1e-11 1e-11 5e-10 1e-09)
VIN_OUTPUT OUTPUT 0 0

* DUT
XU1 INPUT1 INPUT2 OUTPUT NETLIST3

* Loads
CLOAD_INPUT1 INPUT1 0 5e-15

.tran 1e-12 3.0000000000000004e-09
.save time v(INPUT1) v(INPUT2) v(OUTPUT)

.control
  set wr_singlescale
  set filetype=ascii
  run
  wrdata /home/azeem/Desktop/wave-web/wave-backend/run_workspace/runu_ts0b4eks/sim.csv time v(INPUT1) v(INPUT2) v(OUTPUT)
.endc

.end